module ALU;
  
  //Under Progress
endmodule
