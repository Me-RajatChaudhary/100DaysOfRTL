// Code your design here
module day4_alu (
  input logic [7:0]a_i;
  input logic [7:0]b_i;
  input logic [2:0]op;
  output logic [7:0]alu_o
);
  
  
  typedef enum logic
  
  
  
endmodule
