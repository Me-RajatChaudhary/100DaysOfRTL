module 2to1Mux;
