module OddCounter (
);
  
  
  
endmodule
